magic
tech sky130A
timestamp 1628873502
<< nwell >>
rect -120 -52 1957 307
<< ndiff >>
rect 1107 -388 1309 -379
rect 1107 -420 1117 -388
rect 1151 -420 1309 -388
rect 1107 -430 1309 -420
rect 1263 -479 1310 -430
rect 1110 -480 1311 -479
rect 1107 -490 1311 -480
rect 1107 -522 1117 -490
rect 1151 -522 1311 -490
rect 1107 -531 1311 -522
rect 1110 -532 1311 -531
rect -51 -1195 235 -1194
rect -51 -1202 1920 -1195
rect -51 -1205 1710 -1202
rect -51 -1207 712 -1205
rect -51 -1211 90 -1207
rect -51 -1239 -14 -1211
rect 20 -1235 90 -1211
rect 124 -1233 712 -1207
rect 746 -1230 1710 -1205
rect 1744 -1230 1920 -1202
rect 746 -1233 1920 -1230
rect 124 -1235 1920 -1233
rect 20 -1239 1920 -1235
rect -51 -1313 1920 -1239
rect -51 -1315 235 -1313
<< pdiff >>
rect 1758 99 1887 100
rect -78 43 1887 99
rect -78 15 -16 43
rect 16 18 1887 43
rect 16 15 918 18
rect -78 13 918 15
rect -78 -14 94 13
rect 127 11 918 13
rect 127 -14 523 11
rect -78 -17 523 -14
rect -77 -18 523 -17
rect 555 -11 918 11
rect 950 16 1887 18
rect 950 -11 1709 16
rect 555 -13 1709 -11
rect 1741 -13 1887 16
rect 555 -18 1887 -13
rect -77 -25 1887 -18
<< ndiffc >>
rect 1117 -420 1151 -388
rect 1117 -522 1151 -490
rect -14 -1239 20 -1211
rect 90 -1235 124 -1207
rect 712 -1233 746 -1205
rect 1710 -1230 1744 -1202
<< pdiffc >>
rect -16 15 16 43
rect 94 -14 127 13
rect 523 -18 555 11
rect 918 -11 950 18
rect 1709 -13 1741 16
<< poly >>
rect 516 -154 570 -136
rect 78 -174 133 -162
rect 78 -201 91 -174
rect 123 -201 133 -174
rect 78 -336 133 -201
rect 78 -364 86 -336
rect 121 -364 133 -336
rect 516 -182 527 -154
rect 559 -182 570 -154
rect 516 -313 570 -182
rect 516 -341 527 -313
rect 559 -341 570 -313
rect 516 -350 570 -341
rect 904 -146 960 -121
rect 904 -174 917 -146
rect 949 -174 960 -146
rect 904 -310 960 -174
rect 904 -338 917 -310
rect 949 -338 960 -310
rect 904 -349 960 -338
rect 1700 -155 1754 -144
rect 1700 -183 1710 -155
rect 1742 -183 1754 -155
rect 1700 -325 1754 -183
rect 1700 -353 1710 -325
rect 1742 -353 1754 -325
rect 1700 -358 1754 -353
rect 78 -371 133 -364
rect 518 -451 573 -435
rect 518 -479 530 -451
rect 562 -479 573 -451
rect 518 -615 573 -479
rect 518 -643 529 -615
rect 561 -643 573 -615
rect 518 -651 573 -643
rect 911 -454 965 -435
rect 911 -482 923 -454
rect 955 -482 965 -454
rect 911 -614 965 -482
rect 911 -642 922 -614
rect 954 -642 965 -614
rect 911 -650 965 -642
rect 1699 -745 1756 -731
rect 80 -759 142 -747
rect 80 -787 93 -759
rect 125 -787 142 -759
rect 80 -930 142 -787
rect 1699 -773 1711 -745
rect 1743 -773 1756 -745
rect 80 -958 94 -930
rect 128 -958 142 -930
rect 80 -965 142 -958
rect 703 -888 757 -882
rect 703 -916 713 -888
rect 745 -916 757 -888
rect 703 -1060 757 -916
rect 1699 -953 1756 -773
rect 1699 -981 1713 -953
rect 1745 -981 1756 -953
rect 1699 -992 1756 -981
rect 703 -1088 714 -1060
rect 746 -1088 757 -1060
rect 703 -1096 757 -1088
<< polycont >>
rect 91 -201 123 -174
rect 86 -364 121 -336
rect 527 -182 559 -154
rect 527 -341 559 -313
rect 917 -174 949 -146
rect 917 -338 949 -310
rect 1710 -183 1742 -155
rect 1710 -353 1742 -325
rect 530 -479 562 -451
rect 529 -643 561 -615
rect 923 -482 955 -454
rect 922 -642 954 -614
rect 93 -787 125 -759
rect 1711 -773 1743 -745
rect 94 -958 128 -930
rect 713 -916 745 -888
rect 1713 -981 1745 -953
rect 714 -1088 746 -1060
<< locali >>
rect -34 43 26 55
rect -34 15 -16 43
rect 16 15 26 43
rect -34 -1 26 15
rect 85 13 138 20
rect 85 -14 94 13
rect 127 -14 138 13
rect 85 -24 138 -14
rect 515 11 566 22
rect 515 -18 523 11
rect 555 -18 566 11
rect 515 -28 566 -18
rect 908 18 959 28
rect 908 -11 918 18
rect 950 -11 959 18
rect 908 -22 959 -11
rect 1700 16 1751 27
rect 1700 -13 1709 16
rect 1741 -13 1751 16
rect 1700 -23 1751 -13
rect 506 -154 571 -137
rect 60 -174 133 -161
rect 60 -201 91 -174
rect 123 -201 133 -174
rect 506 -182 527 -154
rect 559 -182 571 -154
rect 907 -146 960 -134
rect 907 -174 917 -146
rect 949 -174 960 -146
rect 907 -181 960 -174
rect 1690 -155 1755 -136
rect 506 -194 571 -182
rect 1690 -183 1710 -155
rect 1742 -183 1755 -155
rect 1690 -193 1755 -183
rect 60 -212 133 -201
rect 508 -313 573 -297
rect 73 -336 131 -324
rect 73 -364 86 -336
rect 121 -364 131 -336
rect 508 -341 527 -313
rect 559 -341 573 -313
rect 508 -354 573 -341
rect 897 -310 962 -297
rect 897 -338 917 -310
rect 949 -338 962 -310
rect 897 -354 962 -338
rect 1689 -325 1754 -305
rect 1689 -353 1710 -325
rect 1742 -353 1754 -325
rect 1689 -362 1754 -353
rect 73 -376 131 -364
rect 1108 -388 1160 -379
rect 1108 -420 1117 -388
rect 1151 -420 1160 -388
rect 1108 -429 1160 -420
rect 520 -451 573 -440
rect 520 -479 530 -451
rect 562 -479 573 -451
rect 520 -487 573 -479
rect 911 -454 964 -444
rect 911 -482 923 -454
rect 955 -482 964 -454
rect 911 -491 964 -482
rect 1108 -490 1160 -481
rect 1108 -522 1117 -490
rect 1151 -522 1160 -490
rect 1108 -531 1160 -522
rect 520 -615 571 -605
rect 520 -643 529 -615
rect 561 -643 571 -615
rect 520 -651 571 -643
rect 897 -614 962 -595
rect 897 -642 922 -614
rect 954 -642 962 -614
rect 897 -652 962 -642
rect 1698 -745 1751 -737
rect 75 -759 135 -747
rect 75 -787 93 -759
rect 125 -787 135 -759
rect 1698 -773 1711 -745
rect 1743 -773 1751 -745
rect 1698 -782 1751 -773
rect 75 -797 135 -787
rect 689 -888 754 -871
rect 689 -916 713 -888
rect 745 -916 754 -888
rect 72 -930 139 -919
rect 689 -928 754 -916
rect 72 -958 94 -930
rect 128 -958 139 -930
rect 72 -966 139 -958
rect 1700 -953 1753 -943
rect 1700 -981 1713 -953
rect 1745 -981 1753 -953
rect 1700 -990 1753 -981
rect 690 -1060 755 -1042
rect 690 -1088 714 -1060
rect 746 -1088 755 -1060
rect 690 -1099 755 -1088
rect -25 -1211 28 -1202
rect -25 -1239 -14 -1211
rect 20 -1239 28 -1211
rect -25 -1249 28 -1239
rect 79 -1207 133 -1198
rect 79 -1235 90 -1207
rect 124 -1235 133 -1207
rect 79 -1245 133 -1235
rect 704 -1205 758 -1196
rect 704 -1233 712 -1205
rect 746 -1233 758 -1205
rect 704 -1243 758 -1233
rect 1701 -1202 1755 -1191
rect 1701 -1230 1710 -1202
rect 1744 -1230 1755 -1202
rect 1701 -1238 1755 -1230
<< metal1 >>
rect -73 161 1893 284
rect -52 -3 51 161
rect 1756 160 1884 161
rect 84 24 133 26
rect -50 -29 51 -3
rect 82 20 137 24
rect 82 -55 138 20
rect 80 -127 138 -55
rect 80 -185 137 -127
rect 80 -206 136 -185
rect 513 -194 567 20
rect 906 -23 960 41
rect 905 -133 961 -23
rect 904 -186 962 -133
rect 1699 -189 1753 25
rect 516 -285 570 -256
rect 78 -369 132 -298
rect 78 -373 135 -369
rect 78 -522 136 -373
rect 516 -412 573 -285
rect 517 -440 573 -412
rect 910 -356 966 -278
rect 910 -363 1156 -356
rect 910 -398 1157 -363
rect 517 -493 575 -440
rect 910 -442 966 -398
rect 1108 -420 1157 -398
rect 910 -495 968 -442
rect 1539 -448 1580 -442
rect 1698 -448 1755 -321
rect 1539 -482 1755 -448
rect 79 -791 136 -522
rect 321 -571 566 -520
rect 1108 -536 1157 -488
rect 1539 -502 1581 -482
rect 1540 -536 1581 -502
rect 920 -587 1084 -536
rect 1108 -579 1581 -536
rect 1698 -502 1755 -482
rect 1698 -571 2053 -502
rect 1108 -582 1157 -579
rect 521 -769 578 -596
rect 906 -769 963 -601
rect 1698 -716 1756 -571
rect 1699 -732 1756 -716
rect 519 -814 964 -769
rect 1698 -785 1756 -732
rect 76 -1084 144 -909
rect 701 -921 757 -814
rect 906 -818 963 -814
rect 1703 -967 1754 -934
rect -39 -1480 61 -1194
rect 75 -1248 144 -1084
rect 705 -1246 757 -1045
rect 1703 -1238 1755 -967
rect -50 -1591 1923 -1480
rect -39 -1596 61 -1591
<< labels >>
rlabel metal1 361 -566 379 -527 1 vin1
rlabel metal1 1053 -578 1071 -539 1 vin2
rlabel metal1 1981 -557 1999 -518 1 vout
<< end >>